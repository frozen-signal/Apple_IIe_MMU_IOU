library IEEE;
use IEEE.std_logic_1164.all;

entity MMU_ADDR_DECODER is
    port (
        A     : in std_logic_vector(15 downto 0);
        PHI_0 : in std_logic;

        CXXX_FXXX : out std_logic;
        FXXX_N    : out std_logic;
        EXXX_N    : out std_logic;
        DXXX_N    : out std_logic;
        CXXX      : out std_logic;
        C8_FXX    : out std_logic;
        C8_FXX_N  : out std_logic;
        C0_7XX_N  : out std_logic;
        E_FXXX_N  : out std_logic;
        D_FXXX    : out std_logic;

        -- There is also an address decoder in the IOU. The addresses decoded by
        -- the MMU are prefixed by 'M'. So, MC00X_N is C00X_N, but decoded by the MMU.
        -- The main difference is that the IOU uses the latched address and the MMU uses
        -- the address bus directly.
        MC0XX_N : out std_logic;
        MC3XX   : out std_logic;
        MC00X_N : out std_logic;
        MC01X_N : out std_logic;
        MC04X_N : out std_logic;
        MC05X_N : out std_logic;
        MC06X_N : out std_logic;
        MC07X_N : out std_logic;
        MCFFF_N : out std_logic;

        S_00_1XX    : out std_logic;  -- HIGH when the ADDRESS at the MMU's input is between $0000 - $01FF ($0[0-1]XX)
        S_04_7XX    : out std_logic;  -- HIGH when the ADDRESS at the MMU's input is between $0400 - $07FF ($0[4-7]XX)
        S_2_3XXX    : out std_logic;  -- HIGH when the ADDRESS at the MMU's input is between $2000 - $3FFF ($[2-3]XXX)
        S_01XX_N    : out std_logic
    );
end MMU_ADDR_DECODER;

architecture RTL of MMU_ADDR_DECODER is
    -- S5 stands for Soft 5, a 'soft' 5v. Comes from the Apple II.
    constant S5 : std_logic := '1'; -- Pull-up resistor see MMU_1 @B-4:A4-15

    component LS138 is
        port (
            A, B, C                        : in std_logic;
            G1, G2A_N, G2B_N               : in std_logic;
            Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7 : out std_logic
        );
    end component;

    signal CXXX_FXXX_INT, EXXX_N_INT, E_FXXX_N_INT, FXXX_N_INT, DXXX_N_INT   : std_logic;
    signal CXXX_INT, MC0XX_N_INT, C8_FXX_INT : std_logic;
    signal S_0XXX, S_0XXX_N, S_X1XX, S_X0_1XX, S_X4_7XX : std_logic;
begin
    -- MMU1 @B-4:F4(LS156)
    CXXX_FXXX_INT <= A(15) and A(14);
    FXXX_N_INT    <= not (CXXX_FXXX_INT and A(13) and A(12));
    EXXX_N_INT    <= not (CXXX_FXXX_INT and A(13) and not A(12));
    DXXX_N_INT    <= not (CXXX_FXXX_INT and not A(13) and A(12));
    CXXX_INT      <= CXXX_FXXX_INT and not A(13) and not A(12);
    C8_FXX_INT    <= CXXX_INT and A(11);
    C8_FXX_N      <= not C8_FXX_INT;
    C0_7XX_N      <= not (CXXX_INT and not A(11));

    -- MMU1 @B-34:D4-11 & F3-11
    E_FXXX_N_INT <= FXXX_N_INT and EXXX_N_INT;    -- There seems to be a typo in the schematics: It's labeled E-FXX' but should be E_FXXX'
    D_FXXX       <= E_FXXX_N_INT nand DXXX_N_INT; -- There seems to be a typo in the schematics: It's labeled D-FXXX' (active low) but should be D-FXXX (active high) (see also MMU2 @C-2:D3-9)

    -- MMU1 @C-3:J4
    MC0XX_N_INT <= (not CXXX_INT) or A(11) or (A(10) or A(9) or A(8));
    MC3XX       <= not((not CXXX_INT) or A(11) or (A(10) or (not A(9)) or (not A(8))));

    -- MMU1 @C-3:J5
    MMU_1_J5 : LS138 port map(
        A     => A(4),
        B     => A(5),
        C     => A(6),
        G1    => S5,
        G2A_N => A(7),
        G2B_N => MC0XX_N_INT,
        Y0    => MC00X_N,
        Y1    => MC01X_N,
        Y2    => open,
        Y3    => open,
        Y4    => MC04X_N,
        Y5    => MC05X_N, -- DIFFERENT THAN IN THE EMULATOR SCHEMATICS; Used for the soft switches HIRES (C056/7) and PG2 (C054/5). See the ASIC schematics.
        Y6    => MC06X_N,
        Y7    => MC07X_N
    );

    -- MMU2 @C-4:A2-9
    MCFFF_N <= not (C8_FXX_INT and PHI_0 -- There seems to be a typo in the schematics: Should be C8-FXX instead of C8-FXXX
        and A(10) and A(9) and A(8) and A(7) and A(6)
        and A(5) and A(4) and A(3) and A(2) and A(1) and A(0));

    -- MMU_2 @D-2
    -- Φ0/1XX and Φ0/7XX are only used in the computation of SELMB_N (See MMU_2 @B-1). The computation of SELMB_N in the logical gate schematics seems to have an error.
    -- Using "Apple IIe Diagnostic, v2.1" reports an error while testing AUX RAM. Also, the game "Aliens" will hang while loading. Comparing a logic analyzer trace of the logical schematics vs the official MMU
    -- will reveal a difference on /EN80 and /CASEN.
    -- Instead this implementation will use the ASIC computation of SELMB_N
    -- Also: PHI_0_1XX_N_INT:  There seems to be a typo in the schematics: It's labeled PHI_0_1XX but should be PHI_0_1XX_N (see also MMU2 @C-2:S3-1)

    -- From ASIC Schematics
    S_0XXX <= not (A(15) or A(14) or A(13) or A(12));
    S_0XXX_N <= not S_0XXX;
    S_2_3XXX <= not ((not A(13)) or A(14) or A(15));
    S_X0_1XX <= not (A(11) or A(10) or A(9));
    S_X4_7XX <= not (A(11) or (not A(10)));
    S_X1XX <= not (A(11) or A(10) or A(9) or (not A(8)));

    S_00_1XX <= (not S_X0_1XX) nor S_0XXX_N;
    S_04_7XX <= (not S_X4_7XX) nor S_0XXX_N;
    S_01XX_N <= not (S_0XXX and S_X1XX);

    CXXX_FXXX   <= CXXX_FXXX_INT;
    EXXX_N      <= EXXX_N_INT;
    E_FXXX_N    <= E_FXXX_N_INT;
    FXXX_N      <= FXXX_N_INT;
    DXXX_N      <= DXXX_N_INT;
    CXXX        <= CXXX_INT;
    MC0XX_N     <= MC0XX_N_INT;
    C8_FXX      <= C8_FXX_INT;

end RTL;
